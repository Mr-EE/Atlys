

 
 
 




window new WaveWindow  -name  "Waves for BMG Example Design"
waveform  using  "Waves for BMG Example Design"

      waveform add -signals /bram_tdp_2000d_16wr_8rd_tb/status
      waveform add -signals /bram_tdp_2000d_16wr_8rd_tb/bram_tdp_2000d_16wr_8rd_synth_inst/bmg_port/RSTA
      waveform add -signals /bram_tdp_2000d_16wr_8rd_tb/bram_tdp_2000d_16wr_8rd_synth_inst/bmg_port/CLKA
      waveform add -signals /bram_tdp_2000d_16wr_8rd_tb/bram_tdp_2000d_16wr_8rd_synth_inst/bmg_port/ADDRA
      waveform add -signals /bram_tdp_2000d_16wr_8rd_tb/bram_tdp_2000d_16wr_8rd_synth_inst/bmg_port/DINA
      waveform add -signals /bram_tdp_2000d_16wr_8rd_tb/bram_tdp_2000d_16wr_8rd_synth_inst/bmg_port/WEA
      waveform add -signals /bram_tdp_2000d_16wr_8rd_tb/bram_tdp_2000d_16wr_8rd_synth_inst/bmg_port/ENA
      waveform add -signals /bram_tdp_2000d_16wr_8rd_tb/bram_tdp_2000d_16wr_8rd_synth_inst/bmg_port/DOUTA
      waveform add -signals /bram_tdp_2000d_16wr_8rd_tb/bram_tdp_2000d_16wr_8rd_synth_inst/bmg_port/RSTB
      waveform add -signals /bram_tdp_2000d_16wr_8rd_tb/bram_tdp_2000d_16wr_8rd_synth_inst/bmg_port/CLKB
      waveform add -signals /bram_tdp_2000d_16wr_8rd_tb/bram_tdp_2000d_16wr_8rd_synth_inst/bmg_port/ADDRB
      waveform add -signals /bram_tdp_2000d_16wr_8rd_tb/bram_tdp_2000d_16wr_8rd_synth_inst/bmg_port/ENB
      waveform add -signals /bram_tdp_2000d_16wr_8rd_tb/bram_tdp_2000d_16wr_8rd_synth_inst/bmg_port/DINB
      waveform add -signals /bram_tdp_2000d_16wr_8rd_tb/bram_tdp_2000d_16wr_8rd_synth_inst/bmg_port/WEB
      waveform add -signals /bram_tdp_2000d_16wr_8rd_tb/bram_tdp_2000d_16wr_8rd_synth_inst/bmg_port/DOUTB

console submit -using simulator -wait no "run"
